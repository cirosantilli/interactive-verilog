module main(input in1, input in2, output out);
    wire in1, in2, out;
    assign out = in1 & in2;
endmodule
